----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 20.07.2024 14:56:57
-- Design Name: 
-- Module Name: nueron_sigmoid - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
library work;
use work.utilities.all;
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity nn is
Port ( input : in STD_LOGIC_VECTOR (29 downto 0);          
       led_ans : out STD_LOGIC
       );
end nn;

architecture Behavioral of nn is
signal in_layer2 : std_logic_vector(233 downto 0) := (others => '0');
constant m : matrix(0 to 8) :=(("00000000000000000100001011", "00000000000000000001100000", "00000000000000000011010001", "00000000000000000101000010", "00000000000000000001111101", "00000000000000000011101100", "00000000000000000001001000", "00000000000000000000110010", "00000000000000000010000111", "00000000000000000010111000"),
("00000000000000000000101001", "00000000000000000011000111", "00000000000000000011100100", "00000000000000000011010110", "00000000000000000100101010", "00000000000000000010000000", "00000000000000000010111010", "00000000000000000001010010", "00000000000000000001101101", "00000000000000000010010100"),
("00000000000000000110011000", "00000000000000000011000100", "00000000000000000011110100", "00000000000000000101100111", "00000000000000000100100001", "00000000000000000010010001", "00000000000000000101010001", "00000000000000000011001001", "00000000000000000011100010", "00000000000000000010111001"),
("00000000000000000110000011", "00000000000000000010001101", "00000000000000000001111111", "00000000000000000010000001", "00000000000000000000111010", "00000000000000000000111011", "00000000000000000101011000", "00000000000000000101110111", "00000000000000000010110011", "00000000000000000011100101"),
("00000000000000000110000010", "00000000000000000001001000", "00000000000000000100111111", "00000000000000000010011100", "00000000000000000010100010", "00000000000000000000101110", "00000000000000000011101000", "00000000000000000011110011", "00000000000000000011001001", "00000000000000000010001000"),
("00000000000000000101000100", "00000000000000000011011000", "00000000000000000101010001", "00000000000000000001001101", "00000000000000000001011010", "00000000000000000011100001", "00000000000000000001000000", "00000000000000000000110000", "00000000000000000010000110", "00000000000000000110000010"),
("00000000000000000110000101", "00000000000000000100001011", "00000000000000000001001011", "00000000000000000001111000", "00000000000000000110000111", "00000000000000000001101110", "00000000000000000011111000", "00000000000000000001110011", "00000000000000000100010100", "00000000000000000011100001"),
("00000000000000000010001101", "00000000000000000101101011", "00000000000000000011001000", "00000000000000000010100000", "00000000000000000010011010", "00000000000000000100011101", "00000000000000000011101001", "00000000000000000010011000", "00000000000000000101110101", "00000000000000000010110111"),
("11111111111111001001010010", "11111111111111101111111010", "11111111111111011101101010", "00000000000000101100001101", "00000000000000011010101110", "11111111111111111111001011", "00000000000000100001000110", "00000000000000001111100111", "00000000000000000001011110", "00000000000000000000000000"));

-- 0 to 8 are weights for 1st layer nueron, 9 is the weights for second layer nueron and the last vector in 
-- 9th weight has to be just 0 
signal output: std_logic_vector(25 downto 0) := (others => '0');
begin
layer1_nuer : for i in 0 to 7 generate
      NUERx : entity work.nueron(layer1)
              generic map(w => m(i), in_size => 30)
              port map(input => input, output => in_layer2(i*26 + 25 downto i*26));
              end generate;
-- adding the bias term 
in_layer2(233 downto 208) <= "00000000000001000000000000";
NUER_LAY2 : entity work.nueron(layer2)
            generic map(w => m(8), in_size =>234)
            port map(input=>in_layer2(233 downto 0), output => output);
        
COMPARE : process(output)
          variable threshhold : std_logic_vector(25 downto 0):= "00000000000000100000000000";
          begin
          if unsigned(output) > unsigned(threshhold) then
          led_ans <= '1';
          else
          led_ans <= '0';
          end if;
          end process COMPARE;          
end Behavioral;
